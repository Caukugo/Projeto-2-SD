module Testando (
    input [4:0] a, b,
    output [4:0] f
);

assign f = a & b;


endmodule